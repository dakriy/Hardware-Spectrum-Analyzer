----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:09:45 12/05/2018 
-- Design Name: 
-- Module Name:    ROM - ROM_arch 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

use Spectrum_Analyzer.all;

entity ROM is
	port(
		dataout : out rom_dat_type(0 to 31);
		addr : in std_logic_vector(3 downto 0)
	);
end ROM;

architecture ROM_arch of ROM is
	type rom_type is arraY (0 to 15) of rom_dat_type(0 to 31);
	signal read_only_memory : rom_type :=
	(
		(
			X"2B5",
			X"153",
			X"19D",
			X"1EC",
			X"23D",
			X"290",
			X"2E4",
			X"335",
			X"385",
			X"3CE",
			X"40F",
			X"44A",
			X"47A",
			X"49F",
			X"4B8",
			X"4C5",
			X"4C5",
			X"4B8",
			X"49F",
			X"47A",
			X"44A",
			X"40F",
			X"3CE",
			X"385",
			X"335",
			X"2E4",
			X"290",
			X"23D",
			X"1EC",
			X"19D",
			X"153",
			X"2B5"
		),
		(
			X"177",
			X"F3B",
			X"EC4",
			X"E15",
			X"D55",
			X"CAE",
			X"C4B",
			X"C4F",
			X"CD1",
			X"DD3",
			X"F44",
			X"0FD",
			X"2C9",
			X"46B",
			X"5A8",
			X"653",
			X"653",
			X"5A8",
			X"46B",
			X"2C9",
			X"0FD",
			X"F44",
			X"DD3",
			X"CD1",
			X"C4F",
			X"C4B",
			X"CAE",
			X"D55",
			X"E15",
			X"EC4",
			X"F3B",
			X"177"
		),
		(
			X"02A",
			X"13D",
			X"13A",
			X"171",
			X"12D",
			X"072",
			X"F51",
			X"E07",
			X"CF1",
			X"C6A",
			X"CB6",
			X"DE0",
			X"FB3",
			X"1C4",
			X"38D",
			X"495",
			X"495",
			X"38D",
			X"1C4",
			X"FB3",
			X"DE0",
			X"CB6",
			X"C6A",
			X"CF1",
			X"E07",
			X"F51",
			X"072",
			X"12D",
			X"171",
			X"13A",
			X"13D",
			X"02A"
		),
		(
			X"FB2",
			X"EAF",
			X"F11",
			X"F6C",
			X"084",
			X"1BB",
			X"27B",
			X"22E",
			X"0B5",
			X"E8F",
			X"CB1",
			X"C14",
			X"D30",
			X"FAB",
			X"276",
			X"448",
			X"448",
			X"276",
			X"FAB",
			X"D30",
			X"C14",
			X"CB1",
			X"E8F",
			X"0B5",
			X"22E",
			X"27B",
			X"1BB",
			X"084",
			X"F6C",
			X"F11",
			X"EAF",
			X"FB2"
		),
		(
			X"08D",
			X"144",
			X"05A",
			X"F7D",
			X"E37",
			X"E26",
			X"F80",
			X"1B9",
			X"328",
			X"27D",
			X"FCF",
			X"CDD",
			X"BD8",
			X"DB7",
			X"153",
			X"426",
			X"426",
			X"153",
			X"DB7",
			X"BD8",
			X"CDD",
			X"FCF",
			X"27D",
			X"328",
			X"1B9",
			X"F80",
			X"E26",
			X"E37",
			X"F7D",
			X"05A",
			X"144",
			X"08D"
		),
		(
			X"E68",
			X"E04",
			X"0B6",
			X"29D",
			X"329",
			X"F5D",
			X"B77",
			X"B3A",
			X"093",
			X"64A",
			X"663",
			X"F96",
			X"876",
			X"86E",
			X"027",
			X"7FF",
			X"7FF",
			X"027",
			X"86E",
			X"876",
			X"F96",
			X"663",
			X"64A",
			X"093",
			X"B3A",
			X"B77",
			X"F5D",
			X"329",
			X"29D",
			X"0B6",
			X"E04",
			X"E68"
		),
		(
			X"106",
			X"081",
			X"F19",
			X"E93",
			X"010",
			X"22C",
			X"185",
			X"E6A",
			X"CD0",
			X"FA1",
			X"374",
			X"2F8",
			X"E35",
			X"B86",
			X"EC8",
			X"3D2",
			X"3D2",
			X"EC8",
			X"B86",
			X"E35",
			X"2F8",
			X"374",
			X"FA1",
			X"CD0",
			X"E6A",
			X"185",
			X"22C",
			X"010",
			X"E93",
			X"F19",
			X"081",
			X"106"
		),
		(
			X"F08",
			X"006",
			X"150",
			X"0AF",
			X"E7C",
			X"EA3",
			X"1B7",
			X"285",
			X"ED5",
			X"CA0",
			X"058",
			X"41A",
			X"10C",
			X"BF1",
			X"DAA",
			X"38D",
			X"38D",
			X"DAA",
			X"BF1",
			X"10C",
			X"41A",
			X"058",
			X"CA0",
			X"ED5",
			X"285",
			X"1B7",
			X"EA3",
			X"E7C",
			X"0AF",
			X"150",
			X"006",
			X"F08"
		),
		(
			X"1A1",
			X"EF4",
			X"D61",
			X"0E6",
			X"328",
			X"DFC",
			X"B7C",
			X"2B6",
			X"555",
			X"C2B",
			X"9D4",
			X"4C4",
			X"68E",
			X"A51",
			X"95B",
			X"64D",
			X"64D",
			X"95B",
			X"A51",
			X"68E",
			X"4C4",
			X"9D4",
			X"C2B",
			X"555",
			X"2B6",
			X"B7C",
			X"DFC",
			X"328",
			X"0E6",
			X"D61",
			X"EF4",
			X"1A1"
		),
		(
			X"F5F",
			X"0EE",
			X"0DF",
			X"EBE",
			X"FBC",
			X"224",
			X"F63",
			X"D8E",
			X"201",
			X"20E",
			X"CA7",
			X"F32",
			X"423",
			X"F01",
			X"C0B",
			X"2CA",
			X"2CA",
			X"C0B",
			X"F01",
			X"423",
			X"F32",
			X"CA7",
			X"20E",
			X"201",
			X"D8E",
			X"F63",
			X"224",
			X"FBC",
			X"EBE",
			X"0DF",
			X"0EE",
			X"F5F"
		),
		(
			X"069",
			X"ED1",
			X"FD5",
			X"14A",
			X"EBD",
			X"F40",
			X"263",
			X"ED1",
			X"E04",
			X"330",
			X"F9D",
			X"CA4",
			X"33F",
			X"0FE",
			X"BBA",
			X"269",
			X"269",
			X"BBA",
			X"0FE",
			X"33F",
			X"CA4",
			X"F9D",
			X"330",
			X"E04",
			X"ED1",
			X"263",
			X"F40",
			X"EBD",
			X"14A",
			X"FD5",
			X"ED1",
			X"069"
		),
		(
			X"FD4",
			X"13E",
			X"F74",
			X"F76",
			X"1AB",
			X"E90",
			X"F96",
			X"26D",
			X"D79",
			X"025",
			X"2D6",
			X"C6D",
			X"10C",
			X"2B2",
			X"BC7",
			X"203",
			X"203",
			X"BC7",
			X"2B2",
			X"10C",
			X"C6D",
			X"2D6",
			X"025",
			X"D79",
			X"26D",
			X"F96",
			X"E90",
			X"1AB",
			X"F76",
			X"F74",
			X"13E",
			X"FD4"
		),
		(
			X"FDB",
			X"DC7",
			X"208",
			X"EFA",
			X"EBA",
			X"39E",
			X"BCF",
			X"1F7",
			X"23B",
			X"A1A",
			X"663",
			X"D2E",
			X"D03",
			X"77D",
			X"852",
			X"339",
			X"339",
			X"852",
			X"77D",
			X"D03",
			X"D2E",
			X"663",
			X"A1A",
			X"23B",
			X"1F7",
			X"BCF",
			X"39E",
			X"EBA",
			X"EFA",
			X"208",
			X"DC7",
			X"FDB"
		),
		(
			X"09D",
			X"1A6",
			X"DD3",
			X"273",
			X"E3F",
			X"FEE",
			X"28D",
			X"B46",
			X"580",
			X"BCF",
			X"0F2",
			X"331",
			X"95F",
			X"7E9",
			X"9A6",
			X"26D",
			X"26D",
			X"9A6",
			X"7E9",
			X"95F",
			X"331",
			X"0F2",
			X"BCF",
			X"580",
			X"B46",
			X"28D",
			X"FEE",
			X"E3F",
			X"273",
			X"DD3",
			X"1A6",
			X"09D"
		),
		(
			X"F15",
			X"EF7",
			X"1B6",
			X"D69",
			X"34F",
			X"C7A",
			X"2F9",
			X"E6F",
			X"F6C",
			X"31C",
			X"A7E",
			X"738",
			X"839",
			X"6F3",
			X"B33",
			X"1B7",
			X"1B7",
			X"B33",
			X"6F3",
			X"839",
			X"738",
			X"A7E",
			X"31C",
			X"F6C",
			X"E6F",
			X"2F9",
			X"C7A",
			X"34F",
			X"D69",
			X"1B6",
			X"EF7",
			X"F15"
		),
		(
			X"EE6",
			X"103",
			X"E96",
			X"1E9",
			X"D91",
			X"2F3",
			X"C98",
			X"3C5",
			X"C03",
			X"40A",
			X"C1B",
			X"38B",
			X"D00",
			X"248",
			X"E93",
			X"07C",
			X"07C",
			X"E93",
			X"248",
			X"D00",
			X"38B",
			X"C1B",
			X"40A",
			X"C03",
			X"3C5",
			X"C98",
			X"2F3",
			X"D91",
			X"1E9",
			X"E96",
			X"103",
			X"EE6"
		)
);
begin

		dataout <= read_only_memory(to_integer(unsigned(addr)));

end ROM_arch;

